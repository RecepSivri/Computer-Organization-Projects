library verilog;
use verilog.vl_types.all;
entity fullAdder_4bit is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end fullAdder_4bit;
