library verilog;
use verilog.vl_types.all;
entity project4 is
    port(
        a               : in     vl_logic
    );
end project4;
