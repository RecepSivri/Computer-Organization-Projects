library verilog;
use verilog.vl_types.all;
entity substruct_4bit is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end substruct_4bit;
