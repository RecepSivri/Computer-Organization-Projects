library verilog;
use verilog.vl_types.all;
entity demo_main is
end demo_main;
