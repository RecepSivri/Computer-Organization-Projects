library verilog;
use verilog.vl_types.all;
entity mips_core_tester is
    port(
        a               : in     vl_logic
    );
end mips_core_tester;
